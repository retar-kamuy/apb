class apb_base_test extends uvm_test;
  `uvm_component_utils(apb_base_test)

  apb_env env;
  // apb_sequence seq;
  bus_sequence seq;

  function new(string name = "apb_base_test", uvm_component parent=null);
    super.new(name, parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);

    env = apb_env::type_id::create("env", this);
    // seq = apb_sequence::type_id::create("seq");
    seq = bus_sequence::type_id::create("seq");
  endfunction

  task run_phase(uvm_phase phase);
    phase.raise_objection(this);
    seq.start(env.agent.sequencer);
    phase.drop_objection(this);
  endtask

endclass
