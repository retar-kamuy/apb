`ifndef DEFINES_SVH_
`define DEFINES_SVH_

`define ADDR_WIDTH 32
`define DATA_WIDTH 32

`endif  // DEFINES_SVH_
